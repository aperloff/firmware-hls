`timescale 1ns / 1ps

module SectorProcessor(
  input   ap_clk,
  input   ap_rst,
  input   ap_start,
  output   ap_done,
  output   ap_idle,
  output   ap_ready,
  input  [2:0] bx_V,
  output  [7:0] match1_dataarray_data_V_writeaddr,
  output   match1_dataarray_data_V_enb,
  input  [13:0] match1_dataarray_data_V_dout,
  input  [7:0] match1_nentries_0_V,
  input  [7:0] match1_nentries_1_V,
  input  [7:0] match1_nentries_2_V,
  input  [7:0] match1_nentries_3_V,
  input  [7:0] match1_nentries_4_V,
  input  [7:0] match1_nentries_5_V,
  input  [7:0] match1_nentries_6_V,
  input  [7:0] match1_nentries_7_V,
  output  [7:0] match2_dataarray_data_V_writeaddr,
  output   match2_dataarray_data_V_enb,
  input  [13:0] match2_dataarray_data_V_dout,
  input  [7:0] match2_nentries_0_V,
  input  [7:0] match2_nentries_1_V,
  input  [7:0] match2_nentries_2_V,
  input  [7:0] match2_nentries_3_V,
  input  [7:0] match2_nentries_4_V,
  input  [7:0] match2_nentries_5_V,
  input  [7:0] match2_nentries_6_V,
  input  [7:0] match2_nentries_7_V,
  output  [7:0] match3_dataarray_data_V_writeaddr,
  output   match3_dataarray_data_V_enb,
  input  [13:0] match3_dataarray_data_V_dout,
  input  [7:0] match3_nentries_0_V,
  input  [7:0] match3_nentries_1_V,
  input  [7:0] match3_nentries_2_V,
  input  [7:0] match3_nentries_3_V,
  input  [7:0] match3_nentries_4_V,
  input  [7:0] match3_nentries_5_V,
  input  [7:0] match3_nentries_6_V,
  input  [7:0] match3_nentries_7_V,
  output  [7:0] match4_dataarray_data_V_writeaddr,
  output   match4_dataarray_data_V_enb,
  input  [13:0] match4_dataarray_data_V_dout,
  input  [7:0] match4_nentries_0_V,
  input  [7:0] match4_nentries_1_V,
  input  [7:0] match4_nentries_2_V,
  input  [7:0] match4_nentries_3_V,
  input  [7:0] match4_nentries_4_V,
  input  [7:0] match4_nentries_5_V,
  input  [7:0] match4_nentries_6_V,
  input  [7:0] match4_nentries_7_V,
  output  [7:0] match5_dataarray_data_V_writeaddr,
  output   match5_dataarray_data_V_enb,
  input  [13:0] match5_dataarray_data_V_dout,
  input  [7:0] match5_nentries_0_V,
  input  [7:0] match5_nentries_1_V,
  input  [7:0] match5_nentries_2_V,
  input  [7:0] match5_nentries_3_V,
  input  [7:0] match5_nentries_4_V,
  input  [7:0] match5_nentries_5_V,
  input  [7:0] match5_nentries_6_V,
  input  [7:0] match5_nentries_7_V,
  output  [7:0] match6_dataarray_data_V_writeaddr,
  output   match6_dataarray_data_V_enb,
  input  [13:0] match6_dataarray_data_V_dout,
  input  [7:0] match6_nentries_0_V,
  input  [7:0] match6_nentries_1_V,
  input  [7:0] match6_nentries_2_V,
  input  [7:0] match6_nentries_3_V,
  input  [7:0] match6_nentries_4_V,
  input  [7:0] match6_nentries_5_V,
  input  [7:0] match6_nentries_6_V,
  input  [7:0] match6_nentries_7_V,
  output  [7:0] match7_dataarray_data_V_writeaddr,
  output   match7_dataarray_data_V_enb,
  input  [13:0] match7_dataarray_data_V_dout,
  input  [7:0] match7_nentries_0_V,
  input  [7:0] match7_nentries_1_V,
  input  [7:0] match7_nentries_2_V,
  input  [7:0] match7_nentries_3_V,
  input  [7:0] match7_nentries_4_V,
  input  [7:0] match7_nentries_5_V,
  input  [7:0] match7_nentries_6_V,
  input  [7:0] match7_nentries_7_V,
  output  [7:0] match8_dataarray_data_V_writeaddr,
  output   match8_dataarray_data_V_enb,
  input  [13:0] match8_dataarray_data_V_dout,
  input  [7:0] match8_nentries_0_V,
  input  [7:0] match8_nentries_1_V,
  input  [7:0] match8_nentries_2_V,
  input  [7:0] match8_nentries_3_V,
  input  [7:0] match8_nentries_4_V,
  input  [7:0] match8_nentries_5_V,
  input  [7:0] match8_nentries_6_V,
  input  [7:0] match8_nentries_7_V,
  output  [9:0] allstub_dataarray_data_V_writeaddr,
  output   allstub_dataarray_data_V_enb,
  input  [61:0] allstub_dataarray_data_V_dout,
  input  [7:0] allstub_nentries_0_V,
  input  [7:0] allstub_nentries_1_V,
  input  [7:0] allstub_nentries_2_V,
  input  [7:0] allstub_nentries_3_V,
  input  [7:0] allstub_nentries_4_V,
  input  [7:0] allstub_nentries_5_V,
  input  [7:0] allstub_nentries_6_V,
  input  [7:0] allstub_nentries_7_V,
  output  [9:0] allproj_dataarray_data_V_writeaddr,
  output   allproj_dataarray_data_V_enb,
  input  [61:0] allproj_dataarray_data_V_dout,
  input  [7:0] allproj_nentries_0_V,
  input  [7:0] allproj_nentries_1_V,
  input  [7:0] allproj_nentries_2_V,
  input  [7:0] allproj_nentries_3_V,
  input  [7:0] allproj_nentries_4_V,
  input  [7:0] allproj_nentries_5_V,
  input  [7:0] allproj_nentries_6_V,
  input  [7:0] allproj_nentries_7_V,
  input  [2:0] bx_o_V,
  output  [7:0] fullmatch1_dataarray_data_V_writeaddr,
  output   fullmatch1_dataarray_data_V_we0,
  output  [44:0] fullmatch1_dataarray_data_V_din,
  output  [7:0] fullmatch1_nentries_0_V,
  output   fullmatch1_nentries_0_V_ap_vld,
  output  [7:0] fullmatch1_nentries_1_V,
  output   fullmatch1_nentries_1_V_ap_vld,
  output  [7:0] fullmatch1_nentries_2_V,
  output   fullmatch1_nentries_2_V_ap_vld,
  output  [7:0] fullmatch1_nentries_3_V,
  output   fullmatch1_nentries_3_V_ap_vld,
  output  [7:0] fullmatch1_nentries_4_V,
  output   fullmatch1_nentries_4_V_ap_vld,
  output  [7:0] fullmatch1_nentries_5_V,
  output   fullmatch1_nentries_5_V_ap_vld,
  output  [7:0] fullmatch1_nentries_6_V,
  output   fullmatch1_nentries_6_V_ap_vld,
  output  [7:0] fullmatch1_nentries_7_V,
  output   fullmatch1_nentries_7_V_ap_vld,
  output  [7:0] fullmatch2_dataarray_data_V_writeaddr,
  output   fullmatch2_dataarray_data_V_we0,
  output  [44:0] fullmatch2_dataarray_data_V_din,
  output  [7:0] fullmatch2_nentries_0_V,
  output   fullmatch2_nentries_0_V_ap_vld,
  output  [7:0] fullmatch2_nentries_1_V,
  output   fullmatch2_nentries_1_V_ap_vld,
  output  [7:0] fullmatch2_nentries_2_V,
  output   fullmatch2_nentries_2_V_ap_vld,
  output  [7:0] fullmatch2_nentries_3_V,
  output   fullmatch2_nentries_3_V_ap_vld,
  output  [7:0] fullmatch2_nentries_4_V,
  output   fullmatch2_nentries_4_V_ap_vld,
  output  [7:0] fullmatch2_nentries_5_V,
  output   fullmatch2_nentries_5_V_ap_vld,
  output  [7:0] fullmatch2_nentries_6_V,
  output   fullmatch2_nentries_6_V_ap_vld,
  output  [7:0] fullmatch2_nentries_7_V,
  output   fullmatch2_nentries_7_V_ap_vld,
  output  [7:0] fullmatch3_dataarray_data_V_writeaddr,
  output   fullmatch3_dataarray_data_V_we0,
  output  [44:0] fullmatch3_dataarray_data_V_din,
  output  [7:0] fullmatch3_nentries_0_V,
  output   fullmatch3_nentries_0_V_ap_vld,
  output  [7:0] fullmatch3_nentries_1_V,
  output   fullmatch3_nentries_1_V_ap_vld,
  output  [7:0] fullmatch3_nentries_2_V,
  output   fullmatch3_nentries_2_V_ap_vld,
  output  [7:0] fullmatch3_nentries_3_V,
  output   fullmatch3_nentries_3_V_ap_vld,
  output  [7:0] fullmatch3_nentries_4_V,
  output   fullmatch3_nentries_4_V_ap_vld,
  output  [7:0] fullmatch3_nentries_5_V,
  output   fullmatch3_nentries_5_V_ap_vld,
  output  [7:0] fullmatch3_nentries_6_V,
  output   fullmatch3_nentries_6_V_ap_vld,
  output  [7:0] fullmatch3_nentries_7_V,
  output   fullmatch3_nentries_7_V_ap_vld,
  output  [7:0] fullmatch4_dataarray_data_V_writeaddr,
  output   fullmatch4_dataarray_data_V_we0,
  output  [44:0] fullmatch4_dataarray_data_V_din,
  output  [7:0] fullmatch4_nentries_0_V,
  output   fullmatch4_nentries_0_V_ap_vld,
  output  [7:0] fullmatch4_nentries_1_V,
  output   fullmatch4_nentries_1_V_ap_vld,
  output  [7:0] fullmatch4_nentries_2_V,
  output   fullmatch4_nentries_2_V_ap_vld,
  output  [7:0] fullmatch4_nentries_3_V,
  output   fullmatch4_nentries_3_V_ap_vld,
  output  [7:0] fullmatch4_nentries_4_V,
  output   fullmatch4_nentries_4_V_ap_vld,
  output  [7:0] fullmatch4_nentries_5_V,
  output   fullmatch4_nentries_5_V_ap_vld,
  output  [7:0] fullmatch4_nentries_6_V,
  output   fullmatch4_nentries_6_V_ap_vld,
  output  [7:0] fullmatch4_nentries_7_V,
  output   fullmatch4_nentries_7_V_ap_vld,
  output  [7:0] fullmatch5_dataarray_data_V_writeaddr,
  output   fullmatch5_dataarray_data_V_we0,
  output  [44:0] fullmatch5_dataarray_data_V_din,
  output  [7:0] fullmatch5_nentries_0_V,
  output   fullmatch5_nentries_0_V_ap_vld,
  output  [7:0] fullmatch5_nentries_1_V,
  output   fullmatch5_nentries_1_V_ap_vld,
  output  [7:0] fullmatch5_nentries_2_V,
  output   fullmatch5_nentries_2_V_ap_vld,
  output  [7:0] fullmatch5_nentries_3_V,
  output   fullmatch5_nentries_3_V_ap_vld,
  output  [7:0] fullmatch5_nentries_4_V,
  output   fullmatch5_nentries_4_V_ap_vld,
  output  [7:0] fullmatch5_nentries_5_V,
  output   fullmatch5_nentries_5_V_ap_vld,
  output  [7:0] fullmatch5_nentries_6_V,
  output   fullmatch5_nentries_6_V_ap_vld,
  output  [7:0] fullmatch5_nentries_7_V,
  output   fullmatch5_nentries_7_V_ap_vld,
  output  [7:0] fullmatch6_dataarray_data_V_writeaddr,
  output   fullmatch6_dataarray_data_V_we0,
  output  [44:0] fullmatch6_dataarray_data_V_din,
  output  [7:0] fullmatch6_nentries_0_V,
  output   fullmatch6_nentries_0_V_ap_vld,
  output  [7:0] fullmatch6_nentries_1_V,
  output   fullmatch6_nentries_1_V_ap_vld,
  output  [7:0] fullmatch6_nentries_2_V,
  output   fullmatch6_nentries_2_V_ap_vld,
  output  [7:0] fullmatch6_nentries_3_V,
  output   fullmatch6_nentries_3_V_ap_vld,
  output  [7:0] fullmatch6_nentries_4_V,
  output   fullmatch6_nentries_4_V_ap_vld,
  output  [7:0] fullmatch6_nentries_5_V,
  output   fullmatch6_nentries_5_V_ap_vld,
  output  [7:0] fullmatch6_nentries_6_V,
  output   fullmatch6_nentries_6_V_ap_vld,
  output  [7:0] fullmatch6_nentries_7_V,
  output   fullmatch6_nentries_7_V_ap_vld,
  output  [7:0] fullmatch7_dataarray_data_V_writeaddr,
  output   fullmatch7_dataarray_data_V_we0,
  output  [44:0] fullmatch7_dataarray_data_V_din,
  output  [7:0] fullmatch7_nentries_0_V,
  output   fullmatch7_nentries_0_V_ap_vld,
  output  [7:0] fullmatch7_nentries_1_V,
  output   fullmatch7_nentries_1_V_ap_vld,
  output  [7:0] fullmatch7_nentries_2_V,
  output   fullmatch7_nentries_2_V_ap_vld,
  output  [7:0] fullmatch7_nentries_3_V,
  output   fullmatch7_nentries_3_V_ap_vld,
  output  [7:0] fullmatch7_nentries_4_V,
  output   fullmatch7_nentries_4_V_ap_vld,
  output  [7:0] fullmatch7_nentries_5_V,
  output   fullmatch7_nentries_5_V_ap_vld,
  output  [7:0] fullmatch7_nentries_6_V,
  output   fullmatch7_nentries_6_V_ap_vld,
  output  [7:0] fullmatch7_nentries_7_V,
  output   fullmatch7_nentries_7_V_ap_vld
);

MatchCalculatorTop_0 MC(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .bx_V(bx_V),
    .match1_dataarray_data_V_address0(match1_dataarray_data_V_writeaddr),
    .match1_dataarray_data_V_ce0(match1_dataarray_data_V_enb),
    .match1_dataarray_data_V_q0(match1_dataarray_data_V_dout),
    .match1_nentries_0_V(match1_nentries_0_V),
    .match1_nentries_1_V(match1_nentries_1_V),
    //.match1_nentries_2_V(match1_nentries_2_V),
    //.match1_nentries_3_V(match1_nentries_3_V),
    //.match1_nentries_4_V(match1_nentries_4_V),
    //.match1_nentries_5_V(match1_nentries_5_V),
    //.match1_nentries_6_V(match1_nentries_6_V),
    //.match1_nentries_7_V(match1_nentries_7_V),
    .match2_dataarray_data_V_address0(match2_dataarray_data_V_writeaddr),
    .match2_dataarray_data_V_ce0(match2_dataarray_data_V_enb),
    .match2_dataarray_data_V_q0(match2_dataarray_data_V_dout),
    .match2_nentries_0_V(match2_nentries_0_V),
    .match2_nentries_1_V(match2_nentries_1_V),
    //.match2_nentries_2_V(match2_nentries_2_V),
    //.match2_nentries_3_V(match2_nentries_3_V),
    //.match2_nentries_4_V(match2_nentries_4_V),
    //.match2_nentries_5_V(match2_nentries_5_V),
    //.match2_nentries_6_V(match2_nentries_6_V),
    //.match2_nentries_7_V(match2_nentries_7_V),
    .match3_dataarray_data_V_address0(match3_dataarray_data_V_writeaddr),
    .match3_dataarray_data_V_ce0(match3_dataarray_data_V_enb),
    .match3_dataarray_data_V_q0(match3_dataarray_data_V_dout),
    .match3_nentries_0_V(match3_nentries_0_V),
    .match3_nentries_1_V(match3_nentries_1_V),
    //.match3_nentries_2_V(match3_nentries_2_V),
    //.match3_nentries_3_V(match3_nentries_3_V),
    //.match3_nentries_4_V(match3_nentries_4_V),
    //.match3_nentries_5_V(match3_nentries_5_V),
    //.match3_nentries_6_V(match3_nentries_6_V),
    //.match3_nentries_7_V(match3_nentries_7_V),
    .match4_dataarray_data_V_address0(match4_dataarray_data_V_writeaddr),
    .match4_dataarray_data_V_ce0(match4_dataarray_data_V_enb),
    .match4_dataarray_data_V_q0(match4_dataarray_data_V_dout),
    .match4_nentries_0_V(match4_nentries_0_V),
    .match4_nentries_1_V(match4_nentries_1_V),
    //.match4_nentries_2_V(match4_nentries_2_V),
    //.match4_nentries_3_V(match4_nentries_3_V),
    //.match4_nentries_4_V(match4_nentries_4_V),
    //.match4_nentries_5_V(match4_nentries_5_V),
    //.match4_nentries_6_V(match4_nentries_6_V),
    //.match4_nentries_7_V(match4_nentries_7_V),
    .match5_dataarray_data_V_address0(match5_dataarray_data_V_writeaddr),
    .match5_dataarray_data_V_ce0(match5_dataarray_data_V_enb),
    .match5_dataarray_data_V_q0(match5_dataarray_data_V_dout),
    .match5_nentries_0_V(match5_nentries_0_V),
    .match5_nentries_1_V(match5_nentries_1_V),
    //.match5_nentries_2_V(match5_nentries_2_V),
    //.match5_nentries_3_V(match5_nentries_3_V),
    //.match5_nentries_4_V(match5_nentries_4_V),
    //.match5_nentries_5_V(match5_nentries_5_V),
    //.match5_nentries_6_V(match5_nentries_6_V),
    //.match5_nentries_7_V(match5_nentries_7_V),
    .match6_dataarray_data_V_address0(match6_dataarray_data_V_writeaddr),
    .match6_dataarray_data_V_ce0(match6_dataarray_data_V_enb),
    .match6_dataarray_data_V_q0(match6_dataarray_data_V_dout),
    .match6_nentries_0_V(match6_nentries_0_V),
    .match6_nentries_1_V(match6_nentries_1_V),
    //.match6_nentries_2_V(match6_nentries_2_V),
    //.match6_nentries_3_V(match6_nentries_3_V),
    //.match6_nentries_4_V(match6_nentries_4_V),
    //.match6_nentries_5_V(match6_nentries_5_V),
    //.match6_nentries_6_V(match6_nentries_6_V),
    //.match6_nentries_7_V(match6_nentries_7_V),
    .match7_dataarray_data_V_address0(match7_dataarray_data_V_writeaddr),
    .match7_dataarray_data_V_ce0(match7_dataarray_data_V_enb),
    .match7_dataarray_data_V_q0(match7_dataarray_data_V_dout),
    .match7_nentries_0_V(match7_nentries_0_V),
    .match7_nentries_1_V(match7_nentries_1_V),
    //.match7_nentries_2_V(match7_nentries_2_V),
    //.match7_nentries_3_V(match7_nentries_3_V),
    //.match7_nentries_4_V(match7_nentries_4_V),
    //.match7_nentries_5_V(match7_nentries_5_V),
    //.match7_nentries_6_V(match7_nentries_6_V),
    //.match7_nentries_7_V(match7_nentries_7_V),
    .match8_dataarray_data_V_address0(match8_dataarray_data_V_writeaddr),
    .match8_dataarray_data_V_ce0(match8_dataarray_data_V_enb),
    .match8_dataarray_data_V_q0(match8_dataarray_data_V_dout),
    .match8_nentries_0_V(match8_nentries_0_V),
    .match8_nentries_1_V(match8_nentries_1_V),
    //.match8_nentries_2_V(match8_nentries_2_V),
    //.match8_nentries_3_V(match8_nentries_3_V),
    //.match8_nentries_4_V(match8_nentries_4_V),
    //.match8_nentries_5_V(match8_nentries_5_V),
    //.match8_nentries_6_V(match8_nentries_6_V),
    //.match8_nentries_7_V(match8_nentries_7_V),
    .allstub_dataarray_data_V_address0(allstub_dataarray_data_V_writeaddr),
    .allstub_dataarray_data_V_ce0(allstub_dataarray_data_V_enb),
    .allstub_dataarray_data_V_q0(allstub_dataarray_data_V_dout),
    .allstub_nentries_0_V(allstub_nentries_0_V),
    .allstub_nentries_1_V(allstub_nentries_1_V),
    .allstub_nentries_2_V(allstub_nentries_2_V),
    .allstub_nentries_3_V(allstub_nentries_3_V),
    .allstub_nentries_4_V(allstub_nentries_4_V),
    .allstub_nentries_5_V(allstub_nentries_5_V),
    .allstub_nentries_6_V(allstub_nentries_6_V),
    .allstub_nentries_7_V(allstub_nentries_7_V),
    .allproj_dataarray_data_V_address0(allproj_dataarray_data_V_writeaddr),
    .allproj_dataarray_data_V_ce0(allproj_dataarray_data_V_enb),
    .allproj_dataarray_data_V_q0(allproj_dataarray_data_V_dout),
    .allproj_nentries_0_V(allproj_nentries_0_V),
    .allproj_nentries_1_V(allproj_nentries_1_V),
    .allproj_nentries_2_V(allproj_nentries_2_V),
    .allproj_nentries_3_V(allproj_nentries_3_V),
    .allproj_nentries_4_V(allproj_nentries_4_V),
    .allproj_nentries_5_V(allproj_nentries_5_V),
    .allproj_nentries_6_V(allproj_nentries_6_V),
    .allproj_nentries_7_V(allproj_nentries_7_V),
    .bx_o_V(bx_o_V),
    .fullmatch1_dataarray_data_V_address0(fullmatch1_dataarray_data_V_writeaddr),
    .fullmatch1_dataarray_data_V_we0(fullmatch1_dataarray_data_V_we0),
    .fullmatch1_dataarray_data_V_d0(fullmatch1_dataarray_data_V_din),
    .fullmatch1_nentries_0_V(fullmatch1_nentries_0_V),
    .fullmatch1_nentries_0_V_ap_vld(fullmatch1_nentries_0_V_ap_vld),
    .fullmatch1_nentries_1_V(fullmatch1_nentries_1_V),
    .fullmatch1_nentries_1_V_ap_vld(fullmatch1_nentries_1_V_ap_vld),
    //.fullmatch1_nentries_2_V(fullmatch1_nentries_2_V),
    //.fullmatch1_nentries_2_V_ap_vld(fullmatch1_nentries_2_V_ap_vld),
    //.fullmatch1_nentries_3_V(fullmatch1_nentries_3_V),
    //.fullmatch1_nentries_3_V_ap_vld(fullmatch1_nentries_3_V_ap_vld),
    //.fullmatch1_nentries_4_V(fullmatch1_nentries_4_V),
    //.fullmatch1_nentries_4_V_ap_vld(fullmatch1_nentries_4_V_ap_vld),
    //.fullmatch1_nentries_5_V(fullmatch1_nentries_5_V),
    //.fullmatch1_nentries_5_V_ap_vld(fullmatch1_nentries_5_V_ap_vld),
    //.fullmatch1_nentries_6_V(fullmatch1_nentries_6_V),
    //.fullmatch1_nentries_6_V_ap_vld(fullmatch1_nentries_6_V_ap_vld),
    //.fullmatch1_nentries_7_V(fullmatch1_nentries_7_V),
    //.fullmatch1_nentries_7_V_ap_vld(fullmatch1_nentries_7_V_ap_vld),
    .fullmatch2_dataarray_data_V_address0(fullmatch2_dataarray_data_V_writeaddr),
    .fullmatch2_dataarray_data_V_we0(fullmatch2_dataarray_data_V_we0),
    .fullmatch2_dataarray_data_V_d0(fullmatch2_dataarray_data_V_din),
    .fullmatch2_nentries_0_V(fullmatch2_nentries_0_V),
    .fullmatch2_nentries_0_V_ap_vld(fullmatch2_nentries_0_V_ap_vld),
    .fullmatch2_nentries_1_V(fullmatch2_nentries_1_V),
    .fullmatch2_nentries_1_V_ap_vld(fullmatch2_nentries_1_V_ap_vld),
    //.fullmatch2_nentries_2_V(fullmatch2_nentries_2_V),
    //.fullmatch2_nentries_2_V_ap_vld(fullmatch2_nentries_2_V_ap_vld),
    //.fullmatch2_nentries_3_V(fullmatch2_nentries_3_V),
    //.fullmatch2_nentries_3_V_ap_vld(fullmatch2_nentries_3_V_ap_vld),
    //.fullmatch2_nentries_4_V(fullmatch2_nentries_4_V),
    //.fullmatch2_nentries_4_V_ap_vld(fullmatch2_nentries_4_V_ap_vld),
    //.fullmatch2_nentries_5_V(fullmatch2_nentries_5_V),
    //.fullmatch2_nentries_5_V_ap_vld(fullmatch2_nentries_5_V_ap_vld),
    //.fullmatch2_nentries_6_V(fullmatch2_nentries_6_V),
    //.fullmatch2_nentries_6_V_ap_vld(fullmatch2_nentries_6_V_ap_vld),
    //.fullmatch2_nentries_7_V(fullmatch2_nentries_7_V),
    //.fullmatch2_nentries_7_V_ap_vld(fullmatch2_nentries_7_V_ap_vld),
    .fullmatch3_dataarray_data_V_address0(fullmatch3_dataarray_data_V_writeaddr),
    .fullmatch3_dataarray_data_V_we0(fullmatch3_dataarray_data_V_we0),
    .fullmatch3_dataarray_data_V_d0(fullmatch3_dataarray_data_V_din),
    .fullmatch3_nentries_0_V(fullmatch3_nentries_0_V),
    .fullmatch3_nentries_0_V_ap_vld(fullmatch3_nentries_0_V_ap_vld),
    .fullmatch3_nentries_1_V(fullmatch3_nentries_1_V),
    .fullmatch3_nentries_1_V_ap_vld(fullmatch3_nentries_1_V_ap_vld),
    //.fullmatch3_nentries_2_V(fullmatch3_nentries_2_V),
    //.fullmatch3_nentries_2_V_ap_vld(fullmatch3_nentries_2_V_ap_vld),
    //.fullmatch3_nentries_3_V(fullmatch3_nentries_3_V),
    //.fullmatch3_nentries_3_V_ap_vld(fullmatch3_nentries_3_V_ap_vld),
    //.fullmatch3_nentries_4_V(fullmatch3_nentries_4_V),
    //.fullmatch3_nentries_4_V_ap_vld(fullmatch3_nentries_4_V_ap_vld),
    //.fullmatch3_nentries_5_V(fullmatch3_nentries_5_V),
    //.fullmatch3_nentries_5_V_ap_vld(fullmatch3_nentries_5_V_ap_vld),
    //.fullmatch3_nentries_6_V(fullmatch3_nentries_6_V),
    //.fullmatch3_nentries_6_V_ap_vld(fullmatch3_nentries_6_V_ap_vld),
    //.fullmatch3_nentries_7_V(fullmatch3_nentries_7_V),
    //.fullmatch3_nentries_7_V_ap_vld(fullmatch3_nentries_7_V_ap_vld),
    .fullmatch4_dataarray_data_V_address0(fullmatch4_dataarray_data_V_writeaddr),
    .fullmatch4_dataarray_data_V_we0(fullmatch4_dataarray_data_V_we0),
    .fullmatch4_dataarray_data_V_d0(fullmatch4_dataarray_data_V_din),
    .fullmatch4_nentries_0_V(fullmatch4_nentries_0_V),
    .fullmatch4_nentries_0_V_ap_vld(fullmatch4_nentries_0_V_ap_vld),
    .fullmatch4_nentries_1_V(fullmatch4_nentries_1_V),
    .fullmatch4_nentries_1_V_ap_vld(fullmatch4_nentries_1_V_ap_vld),
    //.fullmatch4_nentries_2_V(fullmatch4_nentries_2_V),
    //.fullmatch4_nentries_2_V_ap_vld(fullmatch4_nentries_2_V_ap_vld),
    //.fullmatch4_nentries_3_V(fullmatch4_nentries_3_V),
    //.fullmatch4_nentries_3_V_ap_vld(fullmatch4_nentries_3_V_ap_vld),
    //.fullmatch4_nentries_4_V(fullmatch4_nentries_4_V),
    //.fullmatch4_nentries_4_V_ap_vld(fullmatch4_nentries_4_V_ap_vld),
    //.fullmatch4_nentries_5_V(fullmatch4_nentries_5_V),
    //.fullmatch4_nentries_5_V_ap_vld(fullmatch4_nentries_5_V_ap_vld),
    //.fullmatch4_nentries_6_V(fullmatch4_nentries_6_V),
    //.fullmatch4_nentries_6_V_ap_vld(fullmatch4_nentries_6_V_ap_vld),
    //.fullmatch4_nentries_7_V(fullmatch4_nentries_7_V),
    //.fullmatch4_nentries_7_V_ap_vld(fullmatch4_nentries_7_V_ap_vld),
    .fullmatch5_dataarray_data_V_address0(fullmatch5_dataarray_data_V_writeaddr),
    .fullmatch5_dataarray_data_V_we0(fullmatch5_dataarray_data_V_we0),
    .fullmatch5_dataarray_data_V_d0(fullmatch5_dataarray_data_V_din),
    .fullmatch5_nentries_0_V(fullmatch5_nentries_0_V),
    .fullmatch5_nentries_0_V_ap_vld(fullmatch5_nentries_0_V_ap_vld),
    .fullmatch5_nentries_1_V(fullmatch5_nentries_1_V),
    .fullmatch5_nentries_1_V_ap_vld(fullmatch5_nentries_1_V_ap_vld),
    //.fullmatch5_nentries_2_V(fullmatch5_nentries_2_V),
    //.fullmatch5_nentries_2_V_ap_vld(fullmatch5_nentries_2_V_ap_vld),
    //.fullmatch5_nentries_3_V(fullmatch5_nentries_3_V),
    //.fullmatch5_nentries_3_V_ap_vld(fullmatch5_nentries_3_V_ap_vld),
    //.fullmatch5_nentries_4_V(fullmatch5_nentries_4_V),
    //.fullmatch5_nentries_4_V_ap_vld(fullmatch5_nentries_4_V_ap_vld),
    //.fullmatch5_nentries_5_V(fullmatch5_nentries_5_V),
    //.fullmatch5_nentries_5_V_ap_vld(fullmatch5_nentries_5_V_ap_vld),
    //.fullmatch5_nentries_6_V(fullmatch5_nentries_6_V),
    //.fullmatch5_nentries_6_V_ap_vld(fullmatch5_nentries_6_V_ap_vld),
    //.fullmatch5_nentries_7_V(fullmatch5_nentries_7_V),
    //.fullmatch5_nentries_7_V_ap_vld(fullmatch5_nentries_7_V_ap_vld),
    .fullmatch6_dataarray_data_V_address0(fullmatch6_dataarray_data_V_writeaddr),
    .fullmatch6_dataarray_data_V_we0(fullmatch6_dataarray_data_V_we0),
    .fullmatch6_dataarray_data_V_d0(fullmatch6_dataarray_data_V_din),
    .fullmatch6_nentries_0_V(fullmatch6_nentries_0_V),
    .fullmatch6_nentries_0_V_ap_vld(fullmatch6_nentries_0_V_ap_vld),
    .fullmatch6_nentries_1_V(fullmatch6_nentries_1_V),
    .fullmatch6_nentries_1_V_ap_vld(fullmatch6_nentries_1_V_ap_vld),
    //.fullmatch6_nentries_2_V(fullmatch6_nentries_2_V),
    //.fullmatch6_nentries_2_V_ap_vld(fullmatch6_nentries_2_V_ap_vld),
    //.fullmatch6_nentries_3_V(fullmatch6_nentries_3_V),
    //.fullmatch6_nentries_3_V_ap_vld(fullmatch6_nentries_3_V_ap_vld),
    //.fullmatch6_nentries_4_V(fullmatch6_nentries_4_V),
    //.fullmatch6_nentries_4_V_ap_vld(fullmatch6_nentries_4_V_ap_vld),
    //.fullmatch6_nentries_5_V(fullmatch6_nentries_5_V),
    //.fullmatch6_nentries_5_V_ap_vld(fullmatch6_nentries_5_V_ap_vld),
    //.fullmatch6_nentries_6_V(fullmatch6_nentries_6_V),
    //.fullmatch6_nentries_6_V_ap_vld(fullmatch6_nentries_6_V_ap_vld),
    //.fullmatch6_nentries_7_V(fullmatch6_nentries_7_V),
    //.fullmatch6_nentries_7_V_ap_vld(fullmatch6_nentries_7_V_ap_vld),
    .fullmatch7_dataarray_data_V_address0(fullmatch7_dataarray_data_V_writeaddr),
    .fullmatch7_dataarray_data_V_we0(fullmatch7_dataarray_data_V_we0),
    .fullmatch7_dataarray_data_V_d0(fullmatch7_dataarray_data_V_din),
    .fullmatch7_nentries_0_V(fullmatch7_nentries_0_V),
    .fullmatch7_nentries_0_V_ap_vld(fullmatch7_nentries_0_V_ap_vld),
    .fullmatch7_nentries_1_V(fullmatch7_nentries_1_V),
    .fullmatch7_nentries_1_V_ap_vld(fullmatch7_nentries_1_V_ap_vld)
    //.fullmatch7_nentries_2_V(fullmatch7_nentries_2_V),
    //.fullmatch7_nentries_2_V_ap_vld(fullmatch7_nentries_2_V_ap_vld),
    //.fullmatch7_nentries_3_V(fullmatch7_nentries_3_V),
    //.fullmatch7_nentries_3_V_ap_vld(fullmatch7_nentries_3_V_ap_vld),
    //.fullmatch7_nentries_4_V(fullmatch7_nentries_4_V),
    //.fullmatch7_nentries_4_V_ap_vld(fullmatch7_nentries_4_V_ap_vld),
    //.fullmatch7_nentries_5_V(fullmatch7_nentries_5_V),
    //.fullmatch7_nentries_5_V_ap_vld(fullmatch7_nentries_5_V_ap_vld),
    //.fullmatch7_nentries_6_V(fullmatch7_nentries_6_V),
    //.fullmatch7_nentries_6_V_ap_vld(fullmatch7_nentries_6_V_ap_vld),
    //.fullmatch7_nentries_7_V(fullmatch7_nentries_7_V),
    //.fullmatch7_nentries_7_V_ap_vld(fullmatch7_nentries_7_V_ap_vld)
);

endmodule
